module foo(
    input a,
    b,
    inout c,
    d,
    output e,
    f
);

endmodule