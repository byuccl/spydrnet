module foo(
    input a
);

endmodule