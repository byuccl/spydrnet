module foo(
    a,
    b,
    c,
    d,
    e,
    f
);

input a;
input b;
inout c;
inout d;
output e;
output f;

endmodule